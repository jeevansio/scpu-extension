library verilog;
use verilog.vl_types.all;
entity pcpu_tb is
end pcpu_tb;
